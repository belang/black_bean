`timescale 1ns/1ps
// file name: ir_decoder_ir_addr.v
// author: lianghy
// time: 2017-4-19 11:33:16

module ir_decoder_ir_addr(
input clk,
input rst_n,
);
endmodule
