`timescale 1ns/1ps
// file name: black_bean.v
// author: lianghy
// time: 2017-5-17 10:21:01

`include "define.v"

module black_bean(
clk,
rst_n,
);
input clk, rst_n;

controller controller_0(
);

computer computer_0(
);
endmodule
